module InstructionMemory_str(Address, Instruction);
	input [31:0] Address;
	output reg [31:0] Instruction=0;
	
	always @(*)
		case (Address[9:2])
            8'd0: Instruction <= 32'h24080000;
            8'd1: Instruction <= 32'h24090000;
            8'd2: Instruction <= 32'h240a0000;
            8'd3: Instruction <= 32'h240d0000;
            8'd4: Instruction <= 32'h00057021;
            8'd5: Instruction <= 32'h8dcc0000;
            8'd6: Instruction <= 32'h11800003;
            8'd7: Instruction <= 32'h21ad0001;
            8'd8: Instruction <= 32'h21ce0004;
            8'd9: Instruction <= 32'h08000005;
            8'd10: Instruction <= 32'h000d2021;
            8'd11: Instruction <= 32'h240d0000;
            8'd12: Instruction <= 32'h00077021;
            8'd13: Instruction <= 32'h8dcc0000;
            8'd14: Instruction <= 32'h11800003;
            8'd15: Instruction <= 32'h21ad0001;
            8'd16: Instruction <= 32'h21ce0004;
            8'd17: Instruction <= 32'h0800000d;
            8'd18: Instruction <= 32'h000d3021;
            8'd19: Instruction <= 32'h23bdffdc;
            8'd20: Instruction <= 32'hafab0020;
            8'd21: Instruction <= 32'hafaa001c;
            8'd22: Instruction <= 32'hafa90018;
            8'd23: Instruction <= 32'hafa80014;
            8'd24: Instruction <= 32'hafbf0010;
            8'd25: Instruction <= 32'hafa4000c;
            8'd26: Instruction <= 32'hafa50008;
            8'd27: Instruction <= 32'hafa60004;
            8'd28: Instruction <= 32'hafa70000;
            8'd29: Instruction <= 32'h000b2021;
            8'd30: Instruction <= 32'h00062821;
            8'd31: Instruction <= 32'h00073021;
            8'd32: Instruction <= 32'h0c00004e;
            8'd33: Instruction <= 32'h8fab0020;
            8'd34: Instruction <= 32'h8faa001c;
            8'd35: Instruction <= 32'h8fa90018;
            8'd36: Instruction <= 32'h8fa80014;
            8'd37: Instruction <= 32'h8fbf0010;
            8'd38: Instruction <= 32'h8fa4000c;
            8'd39: Instruction <= 32'h8fa50008;
            8'd40: Instruction <= 32'h8fa60004;
            8'd41: Instruction <= 32'h8fa70000;
            8'd42: Instruction <= 32'h23bd0024;
            8'd43: Instruction <= 32'h0104602a;
            8'd44: Instruction <= 32'h1180001f;
            8'd45: Instruction <= 32'h00096880;
            8'd46: Instruction <= 32'h01a76820;
            8'd47: Instruction <= 32'h8dad0000;
            8'd48: Instruction <= 32'h00087080;
            8'd49: Instruction <= 32'h01c57020;
            8'd50: Instruction <= 32'h8dce0000;
            8'd51: Instruction <= 32'h01ae6822;
            8'd52: Instruction <= 32'h15a0000d;
            8'd53: Instruction <= 32'h01266822;
            8'd54: Instruction <= 32'h21ad0001;
            8'd55: Instruction <= 32'h15a00007;
            8'd56: Instruction <= 32'h214a0001;
            8'd57: Instruction <= 32'h20ceffff;
            8'd58: Instruction <= 32'h000e7080;
            8'd59: Instruction <= 32'h01cb7020;
            8'd60: Instruction <= 32'h8dc90000;
            8'd61: Instruction <= 32'h21080001;
            8'd62: Instruction <= 32'h08000041;
            8'd63: Instruction <= 32'h21080001;
            8'd64: Instruction <= 32'h21290001;
            8'd65: Instruction <= 32'h0800004b;
            8'd66: Instruction <= 32'h00096822;
            8'd67: Instruction <= 32'h01a0682a;
            8'd68: Instruction <= 32'h11a00005;
            8'd69: Instruction <= 32'h212effff;
            8'd70: Instruction <= 32'h000e7080;
            8'd71: Instruction <= 32'h01cb7020;
            8'd72: Instruction <= 32'h8dc90000;
            8'd73: Instruction <= 32'h0800004b;
            8'd74: Instruction <= 32'h21080001;
            8'd75: Instruction <= 32'h0800002b;//////////////
            8'd76: Instruction <= 32'h000a1021;
            8'd77: Instruction <= 32'h08000075;
            8'd78: Instruction <= 32'h24080001;
            8'd79: Instruction <= 32'h24090000;
            8'd80: Instruction <= 32'h10a00022;
            8'd81: Instruction <= 32'h240a0000;
            8'd82: Instruction <= 32'hac8a0000;
            8'd83: Instruction <= 32'h0105502a;
            8'd84: Instruction <= 32'h1140001c;
            8'd85: Instruction <= 32'h00085880;
            8'd86: Instruction <= 32'h01665820;
            8'd87: Instruction <= 32'h8d6b0000;
            8'd88: Instruction <= 32'h00096080;
            8'd89: Instruction <= 32'h01866020;
            8'd90: Instruction <= 32'h8d8c0000;
            8'd91: Instruction <= 32'h016c5822;
            8'd92: Instruction <= 32'h15600007;
            8'd93: Instruction <= 32'h00085880;
            8'd94: Instruction <= 32'h01645820;
            8'd95: Instruction <= 32'h212c0001;
            8'd96: Instruction <= 32'had6c0000;
            8'd97: Instruction <= 32'h21080001;
            8'd98: Instruction <= 32'h21290001;
            8'd99: Instruction <= 32'h08000070;
            8'd100: Instruction <= 32'h00095822;
            8'd101: Instruction <= 32'h0160582a;
            8'd102: Instruction <= 32'h11600005;
            8'd103: Instruction <= 32'h212cffff;
            8'd104: Instruction <= 32'h000c6080;
            8'd105: Instruction <= 32'h01846020;
            8'd106: Instruction <= 32'h8d890000;
            8'd107: Instruction <= 32'h08000070;
            8'd108: Instruction <= 32'h00085880;
            8'd109: Instruction <= 32'h01645820;
            8'd110: Instruction <= 32'had600000;
            8'd111: Instruction <= 32'h21080001;
            8'd112: Instruction <= 32'h08000053;
            8'd113: Instruction <= 32'h24020000;
            8'd114: Instruction <= 32'h03e00008;
            8'd115: Instruction <= 32'h24020001;
            8'd116: Instruction <= 32'h03e00008;
            8'd117: Instruction <= 32'h08000075;
			default: Instruction <= 32'h00000000;
		endcase
		
endmodule
